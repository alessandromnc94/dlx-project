library ieee;
use ieee.std_logic_1164.all;

entity dlx is

end entity dlx;

-- structural architecture
architecture structural of dlx is

begin  -- architecture structural

  component cu_hw is
  end component cu_hw;

  component datapath is
  end component datapath;



end architecture structural;
