LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

<<<<<<< HEAD
USE work.my_arith_functions.ALL;

=======
>>>>>>> b5269eb7a9009e8583aa25f6804745188b2d496f
PACKAGE p4_carries_logic_network_types IS

END PACKAGE;
