LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE mux_n_m_1_types IS
  -- matrix for inputs
  TYPE mux_n_m_1_matrix IS ARRAY (NATURAL RANGE <>) OF STD_LOGIC_VECTOR;

END PACKAGE;
