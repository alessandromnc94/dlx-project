entity exclude_gen is
end entity;

architecture behavioral of exclude_gen is
component rca_n is
end component;
component p4_adder is
end component;
component half_adder is
end component;
component full_adder is
end component;
component alu is
end component;
component comparator is
end component;
component zero_comparator is
end component;
component cu_hw is
end component;
component datapath is
end component;
component divider is
end component;
component dff is
end component;
component and_gate is
end component;
component and_gate_n is
end component;
component and_gate_single_n is
end component;
component or_gate is
end component;
component or_gate_n is
end component;
component or_gate_single_n is
end component;
component xor_gate is
end component;
component xor_gate_n is
end component;
component xor_gate_single_n is
end component;
component nand_gate is
end component;
component nand_gate_n is
end component;
component nand_gate_single_n is
end component;
component nor_gate is
end component;
component nor_gate_n is
end component;
component nor_gate_single_n is
end component;
component xnor_gate is
end component;
component xnor_gate_n is
end component;
component xnor_gate_single_n is
end component;
component not_gate is
end component;
component not_gate_n is
end component;
component logicals is
end component;
component logicals_n is
end component;
component booth_multiplier is
end component;
component mux_n_2_1 is
end component;
component mux_n_4_1 is
end component;
component mux_n_5_1 is
end component;
component mux_n_6_1 is
end component;
component mux_n_8_1 is
end component;
component mux_n_16_1 is
end component;
component pg_network is
end component;
component register_file is
end component;
component register_file_win is
end component;
component register_n is
end component;
component rotator is
end component;
component shifter is
end component;
component sign_extender is
end component;
begin

end architecture;