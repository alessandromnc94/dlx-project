library ieee;
use ieee.std_logic_1164.all;

package booth_generator_types is
  constant shifted_pos : integer := 8;
end package;
