LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

USE work.my_arith_functions.ALL;

PACKAGE p4_carries_logic_network_types IS

END PACKAGE;
