LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE register_file_win_types IS

  TYPE reg_array IS (NATURAL RANGE <>) OF STD_LOGIC_VECTOR;

END PACKAGE;
