LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE booth_generator_types IS
  CONSTANT shifted_pos : INTEGER := 8;
END PACKAGE;
